module mem_align
	(
	input clk, // Clock
 	input rst_n, // Reset
	input [255:0] data_in,
	input [4:0] num_bytes,
	output logic [255:0] data_out
	);
endmodule
