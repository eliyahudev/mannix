module mem_mux_a 
	(
	input clk, // Clock
 	input rst_n, // Reset
	input [15:0][255:0] data_in,
	input data_valid,
	input [18:0] base_addr,
	input last,
	input [3:0] num_of_last_valid,
	output [15:0][255:0] data_out
	);
endmodule
